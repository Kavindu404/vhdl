library verilog;
use verilog.vl_types.all;
entity part2 is
    port(
        Clk             : in     vl_logic;
        S               : in     vl_logic;
        Q               : out    vl_logic
    );
end part2;
