library verilog;
use verilog.vl_types.all;
entity part6_vlg_vec_tst is
end part6_vlg_vec_tst;
