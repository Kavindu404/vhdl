library verilog;
use verilog.vl_types.all;
entity sev_seg_dec_vlg_vec_tst is
end sev_seg_dec_vlg_vec_tst;
